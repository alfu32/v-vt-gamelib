module libgamev

pub fn test_something(){
	println("hello")
}